library verilog;
use verilog.vl_types.all;
entity ParqueaderoUnitario_vlg_vec_tst is
end ParqueaderoUnitario_vlg_vec_tst;
